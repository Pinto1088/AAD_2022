library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity DecoderSerial is

	port(clk   : in std_logic;
		  mIn   : in std_logic_vector(3 downto 0);
		  mOut  : out std_logic;
		  valid : out std_logic);
		  
end DecoderSerial;

begin


architecture Struct of DecoderSerial is


end Struct;